module calculator;
  integer x = 5;
  initial
    $display("%d", x+6);
endmodule